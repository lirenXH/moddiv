`timescale 1ns / 1ns
module  UNS_ADD_256_tb;
  wire [15:0] sum;
  wire carry;  
  reg [15:0] datain;
  reg  clk,rega_we,regb_we,dff_we,clr,regs_we,rega_sel_cyc,regb_sel_cyc,regs_sel_cyc;
  reg [255:0] a,b;
  reg [256:0] correct_sum;
  
  UNS_ADD_256  UNS_ADD_256(sum,carry,datain,clk,rega_we,regb_we,dff_we,clr,regs_we,rega_sel_cyc,regb_sel_cyc,regs_sel_cyc);
  
  //clock generation				   
  initial clk = 1;
  always #50 clk = ~clk;
	
  initial 
    begin 
      #20   a=256'h32C4AE2C_1F198119_5F990446_6A39C994_8FE30BBF_F2660BE1_715A4589_334C74C7;
            b=256'hBC3736A2_F4F6779C_59BDCEE3_6B692153_D0A9877C_C62A4740_02DF32E5_2139F0A0;
            correct_sum=a+b;
            datain=a[15:0];
            rega_we=1'b1;
            rega_sel_cyc=1'b0;
      #100  datain=a[31:16];
      #100  datain=a[47:32];
      #100  datain=a[63:48];
      #100  datain=a[79:64];
      #100  datain=a[95:80];
      #100  datain=a[111:96];
      #100  datain=a[127:112];
      #100  datain=a[143:128];
      #100  datain=a[159:144];
      #100  datain=a[175:160];
      #100  datain=a[191:176];
      #100  datain=a[207:192];
      #100  datain=a[223:208];
      #100  datain=a[239:224];
      #100  datain=a[255:240];      
      #100  rega_we=1'b0;
            regb_we=1'b1;
            regb_sel_cyc=1'b0;
            datain=b[15:0];
      #100  datain=b[31:16];
      #100  datain=b[47:32];
      #100  datain=b[63:48];
      #100  datain=b[79:64];
      #100  datain=b[95:80];
      #100  datain=b[111:96];
      #100  datain=b[127:112];
      #100  datain=b[143:128];
      #100  datain=b[159:144];
      #100  datain=b[175:160];
      #100  datain=b[191:176];
      #100  datain=b[207:192];
      #100  datain=b[223:208];
      #100  datain=b[239:224];
      #100  datain=b[255:240];
      #100  regb_we=1'b0;
            clr=1'b1;            
      #100  clr=1'b0;
            rega_we=1'b1;
            regb_we=1'b1;
            regs_we=1'b1;
            dff_we=1'b1;
            rega_sel_cyc=1'b1;
            regb_sel_cyc=1'b1;
            regs_sel_cyc=1'b0;
      #1600 rega_we=1'b0;
            regb_we=1'b0;
            regs_we=1'b0;
            dff_we=1'b0;
      #100  regs_sel_cyc=1'b1;
            regs_we=1'b1;
      #1600 regs_we=1'b0;
      
      #200  a=256'h8542D69E_4C044F18_E8B92435_BF6FF7DE_45728391_5C45517D_722EDB8B_08F1DFC3;
            b=256'h987968B4_FA32C3FD_2417842E_73BBFEFF_2F3C848B_6831D7E0_EC65228B_3937E498;
            correct_sum=a+b;
            datain=a[15:0];
            rega_we=1'b1;
            rega_sel_cyc=1'b0;
      #100  datain=a[31:16];
      #100  datain=a[47:32];
      #100  datain=a[63:48];
      #100  datain=a[79:64];
      #100  datain=a[95:80];
      #100  datain=a[111:96];
      #100  datain=a[127:112];
      #100  datain=a[143:128];
      #100  datain=a[159:144];
      #100  datain=a[175:160];
      #100  datain=a[191:176];
      #100  datain=a[207:192];
      #100  datain=a[223:208];
      #100  datain=a[239:224];
      #100  datain=a[255:240];      
      #100  rega_we=1'b0;
            regb_we=1'b1;
            regb_sel_cyc=1'b0;
            datain=b[15:0];
      #100  datain=b[31:16];
      #100  datain=b[47:32];
      #100  datain=b[63:48];
      #100  datain=b[79:64];
      #100  datain=b[95:80];
      #100  datain=b[111:96];
      #100  datain=b[127:112];
      #100  datain=b[143:128];
      #100  datain=b[159:144];
      #100  datain=b[175:160];
      #100  datain=b[191:176];
      #100  datain=b[207:192];
      #100  datain=b[223:208];
      #100  datain=b[239:224];
      #100  datain=b[255:240];
      #100  regb_we=1'b0;
            clr=1'b1;            
      #100  clr=1'b0;
            rega_we=1'b1;
            regb_we=1'b1;
            regs_we=1'b1;
            dff_we=1'b1;
            rega_sel_cyc=1'b1;
            regb_sel_cyc=1'b1;
            regs_sel_cyc=1'b0;
      #1600 rega_we=1'b0;
            regb_we=1'b0;
            regs_we=1'b0;
            dff_we=1'b0;
      #100  regs_sel_cyc=1'b1;
            regs_we=1'b1;
      #1600 regs_we=1'b0;      
	    
	    #200  $finish;		
    end					
endmodule 
